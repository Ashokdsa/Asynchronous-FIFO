`ifndef DATA
  `define DATA 8
  `define DEPTH 16
`endif
