`ifndef DATA
  `define DATA 8
  `define RCLK 100
  `define WCLK 100
`endif
